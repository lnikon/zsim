o_1_ 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 

c_0_ 0 1 1 1 1 0 0 1 0 1 0 1 0 0 1 0 

c_1_ 0 1 1 0 0 1 0 1 0 0 1 0 0 0 1 0
