c_0_  0 1 1 0 2 1 3 0 4 1 5 1 6 1 7 0 8 0 9 1 10 1
c_1_  0 0 1 0 2 1 3 1 4 1 5 1 6 0 7 0 8 0 9 1 10 1
